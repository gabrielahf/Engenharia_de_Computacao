library IEEE;
use IEEE.Std_Logic_1164.all;

package p_ula is  
            type op_alu is  
                ( uAND, uOR, uXOR, uSLL, uSRL, uADD, uSUB, uINC, uNEG, uZero, uDEC);
end p_ula;


